`timescale 10ns/10ps
module control_TB();

	reg [31:0] in;
	wire [22:0] out;

	control DUT(
		.in(in),
		.out(out)
	);

	initial begin
		in = 32'b0;
	
		#10 in = 32'b000101_10111_00000_0000_1100_0000_0000; //LW
		#10 in = 32'b000110_10111_00110_0000_1111_1111_1111; //SW
		#10 in = 32'b000100_00010_00011_00101_01010_100000;   //ADD
		#10 in = 32'b000100_00100_00101_00110_01010_100010;  //SUB
		#10 in = 32'b000100_00000_00001_00100_01010_110010;  //MUL
		#10 in = 32'b000100_11000_11000_11000_01010_100100;  //AND
		#10 in = 32'b000100_11000_11000_11000_01010_100101;  //OR
		#10 $stop;
		
	end
endmodule