`timescale 1ns/100ps
module ADDRDecoding_TB();

	wire cs;
	reg [31:0] addr;
	integer i;
	
	ADDRDecoding DUT(
		.cs(cs),
		.addr(addr)
	);
	
	initial
	begin
		for(i = 0; i <= 32'h2FFF; i = i + 1)
		#20 addr = i;				
	end
	
endmodule 